module geraPreset(Us,Ua,T,unid_preset,dez_preset);
	input Us,Ua,T;
	output [3:0]unid_preset;
	output [1:0]dez_preset;
endmodule